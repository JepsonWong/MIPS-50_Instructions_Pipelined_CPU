module ALU(ALUctr,A,B,C,Zero);
  input [4:0] ALUctr;
  input [31:0] A,B;
  output [31:0] C;
  output [2:0] Zero;
  
  reg [31:0] D;
  reg M;
  wire [63:0] A_E,B_E;
  
  assign C=D; 
  assign Zero[0]=(D==32'b0)?1:0;
  assign Zero[1]=(ALUctr==5'b10000)? ((M==1'b0)?1:0):(((D[31]==1'b0)&(D!=32'b0))?1:0);
  assign Zero[2]=(ALUctr==5'b10000)? ((M==1'b1)?1:0):(((D[31]==1'b1)&(D!=32'b0))?1:0);
  assign A_E=(A[31]==1'b0)? ({32'b0,A}):({32'b11111111111111111111111111111111,A});
  assign B_E=(B[31]==1'b0)? {32'b0,B}:{32'b11111111111111111111111111111111,B}; 
     
  always @ (ALUctr or A or B)
  begin
  case(ALUctr)
  5'b00000:D<=A+B;
  5'b00001:D<=A+B;
  5'b00010:D<=A-B;
  5'b00011:D<=A-B;
  5'b00100:D<=A&B;
  5'b00101:D<=A|B;
  5'b00110:D<=A^B;
  5'b00111:D<=~(A|B);
  5'b01000:D<={B[15:0],16'b0};
  5'b01001://begin
  //D=A;
  //for(i=0;i<B[10:6];i=i+1)
  //D=D<<1;
  //end 
  D<=A<<B[10:6];                 
  5'b01010:
 // begin
    //D=A;
    //for(i=0;i<B[10:6];i=i+1)
    //D=D>>1;
  //end 
  D<=A>>B[10:6];          
  5'b01011:
  //begin
    //D=A;
   // for(i=0;i<B[10:6];i=i+1)
    //begin
    //D=D>>1;
    //D[31]=A[31];
  //end
  //end  
  D<=A_E>>B[10:6];
  5'b01100:
  //begin
   // D=B;
  //for(i=0;i<A;i=i+1)
 // begin
  //  D=D<<1;
 // end
 // end
 D<=B<<A;
  5'b01101:
  //begin
  //D=B;
//  for(i=0;i<A;i=i+1)
 // begin
//    D=D>>1;
//  end 
 // end
 D<=B>>A;
  5'b01110:
  //begin
   // D=B;
 // for(i=0;i<A;i=i+1)
  //begin
  //  D=D>>1;
    //D[31]=B[31];
 // end 
  //end 
  D<=B_E>>A;
  5'b01111:D<=A;                    //{{B{A[32]}},A[32:32'd32-B]};
  5'b10000:{M,D}<={1'b0,A}-{1'b0,B};
  default: D<=32'b0;
endcase
end

endmodule 